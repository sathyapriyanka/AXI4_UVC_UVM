





   
           



 